`define FPGA
// `define PROBE

