`define FPGA
`define PROBE

