`define FPGA
`define PROBE

`undef SOPHON_SOFT_RST
