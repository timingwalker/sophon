`define FPGA
`define PROBE
