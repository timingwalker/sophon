`define FPGA
//`define PROBE

